LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.numeric_std.all;

ENTITY status_reg IS
	PORT (
        -- Inputs
        -- Outputs
	);
END ENTITY;

ARCHITECTURE status_reg OF stack IS

BEGIN
END status_reg;
