LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.numeric_std.all;

ENTITY fsr_reg IS
	PORT (
        -- Inputs
        -- Outputs
	);
END ENTITY;

ARCHITECTURE fsr_reg OF fsr_reg IS

BEGIN
END fsr_reg;
