LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.numeric_std.all;

ENTITY pc_reg IS
	PORT (
        -- Inputs
        -- Outputs
	);
END ENTITY;

ARCHITECTURE pc_reg OF pc_reg IS

BEGIN
END pc_reg;
