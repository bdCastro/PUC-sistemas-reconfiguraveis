LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.numeric_std.all;

ENTITY stack IS
	PORT (
        -- Inputs
        -- Outputs
	);
END ENTITY;

ARCHITECTURE stack OF stack IS

BEGIN
END stack;
